*
*
*
*                       LINUX           Tue Apr 12 21:19:14 2016
*
*
*
*  PROGRAM  advgen
*
*  Name           : advgen - Quantus QRC - (64-bit)
*  Version        : 14.2.3-s099
*  Build Date     : Wed Jun 17 00:01:02 PDT 2015
*
*  HSPICE LIBRARY
*
*
*

*
.SUBCKT inverter VSS VDD OUTP INP
*
*
*  caps2d version: 10
*
*
*       TRANSISTOR CARDS
*
*
MI1	OUTP#9	INP#9	VSS#1	VSS#2	nmos_hs_top
MM0	OUTP#1	INP#8	VDD#1	VDD	pmos_hs
*
*
*       RESISTOR AND CAP/DIODE CARDS
*
Rn1	INP#8	INP	   82.3333
Rm2	INP	INP#5	    3.5000
Rm3	OUTP	OUTP#2	    0.4434
Rm4	OUTP#2	OUTP#3	    1.8050
Rm5	OUTP#1	OUTP#2	    3.3333
Rm6	VDD	VDD#1	    4.7506
Rl1	INP#6	INP#5	    3.5000
Rl2	OUTP#3	OUTP#4	    1.7500
Rk1	INP#1	INP#6	    3.5000
Rk2	OUTP#4	OUTP#5	    1.7500
Rj2	OUTP#5	OUTP#6	    1.7500
Ri1	INP#1	INP#2	   12.6800
Ri2	OUTP#7	OUTP#6	    4.5900
Rh1	VSS#1	VSS#3	  525.0000
Rh2	VSS#3	VSS#4	    5.0000
Rh3	VSS#2	VSS#3	   10.0000
Rh4	OUTP#7	OUTP#9	  530.0000
Rg1	INP#9	INP#3	   59.0000
Rf1	INP#3	INP#2	   10.0000
Rf3	VSS	VSS#4	    0.4770
*
*       CAPACITOR CARDS
*
*
C1	VDD	INP#8	6.11163E-17
C2	VDD	INP#9	3.99001E-18
C3	VDD	OUTP#5	3.19681E-17
C4	VDD	OUTP#4	3.2727E-17
C5	VDD	INP#6	3.47146E-17
C6	VDD	OUTP#3	1.41497E-16
C7	VDD	INP#2	1.7151E-17
C8	VDD	INP#3	3.47725E-18
C9	VDD	VSS#4	2.14267E-17
C10	VDD	OUTP#1	2.40316E-18
C11	OUTP#9	VSS#1	1.88234E-18
C12	OUTP#9	INP#9	5.4073E-17
C13	VSS#1	INP#9	6.61547E-17
C14	INP#8	OUTP#3	1.10117E-16
C15	OUTP#9	INP#2	4.11761E-18
C16	OUTP#9	INP#3	1.06464E-17
C17	INP#8	OUTP#1	1.23136E-16
C18	VSS#1	INP#2	4.9911E-18
C19	INP#8	VDD#1	2.42189E-16
C20	OUTP#9	VSS#4	2.13401E-18
C21	VSS#1	INP#3	1.24304E-17
C22	OUTP#5	INP#6	2.37229E-18
C23	OUTP#4	INP#6	1.18786E-17
C24	INP#9	VSS#4	9.94863E-17
C25	OUTP#5	INP#2	2.22423E-18
C26	INP#6	OUTP#3	4.22336E-17
C27	OUTP#5	VSS#4	4.09097E-18
C28	OUTP#5	VDD#1	1.99935E-18
C29	OUTP#4	VSS#4	2.113E-18
C30	INP#6	VSS#4	1.18801E-18
C31	OUTP#4	VDD#1	6.01258E-18
C32	OUTP#3	VSS#4	1.70974E-18
C33	INP#6	VDD#1	1.58327E-17
C34	OUTP#3	VDD#1	1.84589E-16
C35	INP#2	VSS#4	6.33457E-17
C36	INP#3	VSS#4	1.339E-17
C37	VSS#4	VDD#1	1.34019E-18
C38	INP#1	OUTP#7	6.7904E-17
C39	VDD	INP#1	7.10379E-17
C40	INP#6	OUTP#7	2.2109E-18
C41	INP#1	OUTP#3	1.17545E-17
C42	OUTP#7	INP#2	8.12647E-17
C43	VSS#1	OUTP#7	8.9511E-18
C44	VDD	INP	1.0963E-16
C45	OUTP#7	INP#3	1.19874E-17
C46	INP	OUTP#3	5.20202E-17
C47	INP#1	VDD#1	5.79534E-18
C48	OUTP#7	VSS#4	1.91952E-16
C49	INP	OUTP#1	4.15628E-17
C50	VSS#1	INP#1	9.82847E-19
C51	OUTP#7	VDD#1	1.88828E-18
C52	INP#1	OUTP#4	4.59273E-17
C53	VDD	OUTP#7	4.26839E-17
C54	INP	VDD#1	9.63657E-17
C55	INP#1	VSS#4	1.62687E-17
C56	INP#1	OUTP#5	5.58033E-17
C57	INP#9	OUTP#7	1.35577E-16
C58	VDD	VSS#1	4.24411E-19
C59	INP	VSS#4	4.52851E-19
C60	INP#9	OUTP#4	4.07981E-19
C61	OUTP#9	INP#1	6.63208E-19
C62	INP	OUTP#5	8.71578E-19
C63	INP#9	OUTP#5	8.96617E-19
C64	INP	OUTP#7	9.53426E-19
C65	OUTP#3	INP#2	1.09032E-18
C66	OUTP#4	INP#2	1.25832E-18
C67	INP	OUTP#4	1.5059E-18
C68	VDD	VSS	1.43621E-16
C69	INP	VSS	4.19217E-18
C70	INP#8	VSS	2.24804E-18
C71	OUTP#9	VSS	1.71133E-19
C72	INP#9	VSS	1.39605E-17
C73	INP#1	VSS	5.78732E-17
C74	OUTP#5	VSS	2.02189E-17
C75	OUTP#4	VSS	2.09976E-17
C76	INP#6	VSS	1.66009E-17
C77	OUTP#3	VSS	1.99904E-17
C78	OUTP#7	VSS	1.20173E-16
C79	INP#2	VSS	4.6934E-17
C80	INP#3	VSS	1.36241E-18
C81	OUTP#1	VSS	1.53072E-18
C82	VDD#1	VSS	1.80938E-17
*
*
.ENDS inverter
*
