*
*
*
*                       LINUX           Sat Mar 19 17:32:16 2016
*
*
*
*  PROGRAM  advgen
*
*  Name           : advgen - Quantus QRC - (64-bit)
*  Version        : 14.2.3-s099
*  Build Date     : Wed Jun 17 00:01:02 PDT 2015
*
*  HSPICE LIBRARY
*
*
*

*
.SUBCKT S3D_inv OUT VSS VDD IN
*
*
*  caps2d version: 10
*
*
*       TRANSISTOR CARDS
*
*
MX15/M0	VSS#3	IN#8	OUT#9	VSS#4	nmos_hs_top
MM0	OUT#1	IN#10	VDD#6	VDD#5	pmos_hs
*
*
*       RESISTOR AND CAP/DIODE CARDS
*
Rm1	IN#10	IN#11	   30.6750	$L=0.46U	$W=0.15U
Rm2	IN#11	IN#6	    6.2408	$L=0.1495U	$W=0.3U
Rl1	IN#6	IN#7	   10.3693	$L=0.4U	$W=0.26U
Rl2	IN#7	IN#5	7.658E-02	$L=0.1495U	$W=0.64U
Rl3	VDD#6	VDD#5	   10.7123	$L=0.96U	$W=0.32U
Rl5	OUT#1	OUT#2	   10.4576	$L=0.61U	$W=0.32U
Rl6	OUT#2	OUT#3	    3.5702	$L=0.1495U	$W=0.64U
Rk1	VDD#4	VDD#5	    3.5000	$L=0.001U	$W=0.3U
Rk2	IN#5	IN#4	    3.5000	$L=0.001U	$W=0.3U
Rk3	OUT#4	OUT#3	    3.5000	$L=0.001U	$W=0.3U
Rj1	VDD#2	VDD#4	    3.5000	$L=0.001U	$W=0.3U
Rj2	IN#4	IN#1	    3.5000	$L=0.001U	$W=0.3U
Rj3	OUT#5	OUT#4	    3.5000	$L=0.001U	$W=0.3U
Ri1	VDD#1	VDD#2	    7.0000	$L=0.001U	$W=0.3U
Ri2	IN#1	IN#2	    7.0000	$L=0.001U	$W=0.3U
Ri3	OUT#6	OUT#5	    3.5000	$L=0.001U	$W=0.3U
Rh1	VDD#1	VDD#3	    9.1800	$L=0.001U	$W=0.3U
Rh2	IN#3	IN#2	    9.1800	$L=0.001U	$W=0.3U
Rh3	OUT#6	OUT	    9.1800	$L=0.001U	$W=0.3U
Rg1	VSS#3	VSS#1	   70.8750	$L=0.21U	$W=0.32U
Rg3	VSS#4	VSS#1	   10.0000	$L=0.001U	$W=0.32U
Rg4	OUT#8	OUT#9	   80.8750	$L=0.21U	$W=0.32U
Rf1	VSS#1	VSS#2	   10.1925	$L=0.56U	$W=0.32U
Rf2	VSS#2	VSS	2.187E-02	$L=0.149U	$W=1.27U
Rf3	IN#8	IN#9	   10.1650	$L=0.39U	$W=0.26U
Rf4	IN#9	IN#3	3.330E-02	$L=0.1595U	$W=0.78U
Rf5	IN#3	IN	4.231E-03	$L=0.03U	$W=0.78U
Rf6	VDD	VDD#3	    0.1205	$L=0.3505U	$W=0.32U
Rf7	OUT#8	OUT#10	    0.2097	$L=0.61U	$W=0.32U
Rf8	OUT#10	OUT	3.218E-02	$L=0.1495U	$W=0.64U
*
*       CAPACITOR CARDS
*
*
C1	OUT	VDD	1.60153E-17
C2	OUT	IN	1.85064E-17
C3	VDD	IN	1.90086E-18
C4	OUT	VSS#3	5.16963E-19
C5	OUT	VDD#1	8.43483E-18
C6	OUT	IN#1	2.61768E-18
C7	OUT	IN#5	1.42738E-18
C8	VDD	OUT#6	3.10285E-18
C9	IN	OUT#9	1.24932E-18
C10	OUT	IN#3	6.29527E-18
C11	IN	VSS#3	1.24535E-18
C12	OUT	VDD#3	1.10296E-17
C13	IN	OUT#6	9.69755E-18
C14	OUT	VSS#1	4.9687E-18
C15	OUT	IN#8	4.29778E-18
C16	IN	VDD#1	4.78367E-18
C17	OUT	VSS#2	7.92781E-19
C18	IN	OUT#5	1.83589E-18
C19	OUT	IN#9	2.16994E-18
C20	IN	VDD#2	1.58656E-18
C21	IN	OUT#4	1.6311E-18
C22	OUT#9	VSS#3	6.52801E-18
C23	IN	VDD#4	1.58171E-18
C24	VDD	OUT#8	1.32695E-17
C25	VSS#3	OUT#6	5.47166E-19
C26	VDD	VSS#1	4.62509E-18
C27	IN	VDD#3	4.09106E-18
C28	VSS#3	VDD#1	9.60834E-19
C29	IN	OUT#8	1.59015E-17
C30	VDD	VSS#2	9.55102E-19
C31	IN	VSS#1	1.61917E-17
C32	OUT#6	VDD#1	3.39417E-17
C33	VDD	OUT#10	4.63879E-18
C34	OUT#6	IN#1	1.80595E-17
C35	IN	VSS#2	5.69222E-18
C36	OUT#6	VDD#2	7.968E-18
C37	VDD#1	OUT#5	8.67437E-18
C38	VDD#1	IN#1	7.7635E-18
C39	OUT#6	IN#4	8.28794E-18
C40	IN	OUT#10	3.21494E-18
C41	OUT#6	VDD#4	2.6453E-18
C42	OUT#5	IN#1	6.55326E-18
C43	VDD#1	OUT#4	2.82122E-18
C44	OUT#5	VDD#2	1.08088E-17
C45	OUT#9	VDD#3	1.107E-18
C46	OUT#6	IN#5	4.21295E-18
C47	VDD#1	IN#4	4.57337E-18
C48	IN#1	VDD#2	3.24656E-18
C49	VSS#3	IN#3	6.71885E-19
C50	IN#10	OUT#1	1.20905E-16
C51	VSS#3	VDD#3	1.1073E-18
C52	OUT#5	IN#4	1.17132E-17
C53	OUT#9	VSS#1	5.43866E-18
C54	IN#1	OUT#4	2.06978E-18
C55	IN#10	VDD#6	1.24474E-16
C56	OUT#6	IN#3	1.79024E-17
C57	OUT#5	VDD#4	5.82675E-18
C58	VSS#3	OUT#8	4.99757E-18
C59	VDD#2	OUT#4	5.43492E-18
C60	VDD#1	IN#5	3.1435E-18
C61	OUT#6	VDD#3	7.96119E-18
C62	IN#1	VDD#4	1.52956E-18
C63	VDD#2	IN#4	4.20007E-18
C64	OUT#5	IN#5	7.4794E-18
C65	OUT#4	IN#4	5.7561E-18
C66	OUT#6	VSS#1	3.42798E-18
C67	VDD#1	IN#3	7.21838E-18
C68	OUT#4	VDD#4	8.41588E-18
C69	VDD#2	IN#5	3.06364E-18
C70	OUT#5	IN#3	2.48108E-18
C71	IN#4	VDD#4	2.52789E-18
C72	VDD#1	OUT#8	5.26549E-18
C73	OUT#4	IN#5	1.23657E-17
C74	OUT#5	IN#6	1.21231E-18
C75	VDD#1	VSS#1	7.26955E-18
C76	OUT#6	VSS#2	4.19218E-19
C77	IN#1	VDD#3	1.87207E-18
C78	VDD#4	OUT#3	1.32174E-18
C79	VDD#2	IN#3	1.61879E-18
C80	OUT#5	VSS#1	4.55459E-19
C81	VDD#4	IN#5	3.25168E-18
C82	IN#1	OUT#8	1.1231E-18
C83	OUT#3	IN#5	4.9902E-18
C84	IN#1	VSS#1	1.85299E-18
C85	OUT#4	IN#6	3.55592E-18
C86	VDD#1	VSS#2	7.76131E-19
C87	VDD#2	VSS#1	7.03073E-19
C88	OUT#5	VDD#6	1.38206E-18
C89	OUT#4	VSS#1	2.64247E-19
C90	VDD#4	IN#6	1.27287E-18
C91	VDD#2	OUT#1	1.30647E-18
C92	IN#4	VSS#1	5.98372E-19
C93	IN#1	VSS#2	2.86265E-19
C94	OUT#3	IN#6	3.56598E-18
C95	VDD#4	VSS#1	2.6825E-19
C96	OUT#4	VDD#6	2.64967E-18
C97	IN#4	OUT#1	1.18956E-18
C98	IN#4	VDD#6	2.38214E-18
C99	IN#5	VSS#1	4.70791E-19
C100	VDD#4	OUT#1	5.10716E-18
C101	IN#3	VDD#3	2.69941E-18
C102	IN#3	OUT#8	4.17771E-18
C103	IN#5	OUT#1	6.24964E-18
C104	IN#3	VSS#1	5.0231E-18
C105	IN#5	VDD#6	9.54412E-18
C106	VDD#3	OUT#8	1.97842E-17
C107	VDD#3	VSS#1	2.91742E-17
C108	VDD#3	IN#8	1.22304E-18
C109	OUT#8	VSS#1	6.16627E-17
C110	OUT#8	IN#8	2.73997E-17
C111	IN#6	OUT#1	3.33545E-17
C112	VSS#1	IN#8	2.82273E-17
C113	IN#3	VSS#2	5.56092E-19
C114	IN#5	OUT#2	2.27294E-18
C115	IN#6	VDD#6	3.49157E-17
C116	VDD#3	VSS#2	1.25055E-17
C117	OUT#8	VSS#2	2.13495E-18
C118	IN#8	VSS#2	4.31802E-18
C119	OUT#1	VDD#6	5.35706E-17
C120	OUT#8	IN#9	3.25951E-18
C121	VDD#3	OUT#10	1.77683E-18
C122	IN#6	OUT#2	3.12885E-18
C123	VSS#1	IN#9	3.10817E-18
C124	OUT#1	IN#7	1.67688E-18
C125	VSS#1	OUT#10	8.929E-19
C126	VDD#6	IN#7	1.97539E-18
C127	IN#8	OUT#10	2.2662E-18
C128	OUT#1	IN#11	2.10893E-17
C129	VDD#6	IN#11	2.01185E-17
C130	VSS#2	IN#9	2.23297E-18
C131	VSS#2	OUT#10	2.7778E-19
C132	VDD#5	OUT#2	4.73316E-18
C133	IN#6	VDD#5	1.81741E-18
C134	VSS#1	VDD#5	2.5026E-19
C135	VDD#5	OUT#1	2.21987E-17
C136	IN#4	VDD#5	1.29837E-18
C137	IN#5	VDD#5	2.48047E-18
C138	IN#10	VDD#5	1.1728E-17
C139	OUT#6	VDD#5	2.55996E-18
C140	OUT#5	VDD#5	3.40619E-18
C141	OUT#4	VDD#5	8.27615E-18
C142	OUT#3	VDD#5	8.59706E-18
C143	OUT#3	VSS#1	7.17447E-20
C144	OUT#5	VSS#2	8.60298E-20
C145	OUT#9	VSS#2	1.41844E-19
C146	VSS#1	OUT#1	1.56587E-19
C147	OUT#3	VDD#3	1.86163E-19
C148	OUT#8	VDD#5	2.02659E-19
C149	VDD#4	OUT#8	2.05649E-19
C150	VDD#1	OUT#2	2.12413E-19
C151	OUT	VDD#6	2.46171E-19
C152	VDD#2	OUT#2	2.97986E-19
C153	VDD	OUT#4	2.98074E-19
C154	VDD#2	OUT#8	4.13374E-19
C155	VDD#1	OUT#10	4.51743E-19
C156	VDD	OUT#5	5.34506E-19
C157	OUT#4	VDD#3	5.6292E-19
C158	OUT#3	VDD#6	6.29417E-19
C159	VDD#1	OUT#1	6.68615E-19
C160	VDD#2	OUT#3	7.24026E-19
C161	OUT	VDD#4	8.33186E-19
C162	OUT#6	VDD#6	8.45715E-19
C163	VDD#4	OUT#2	8.79717E-19
C164	OUT#5	VDD#3	9.65086E-19
C165	OUT#9	VDD#1	9.75592E-19
C166	OUT	VDD#2	9.97344E-19
C167	VDD#1	OUT#3	1.00526E-18
C168	OUT	VDD#5	1.07418E-18
C169	IN#4	OUT#10	9.02231E-20
C170	IN#5	OUT#10	1.12077E-19
C171	OUT#6	IN#7	1.2017E-19
C172	IN	OUT#3	1.34913E-19
C173	OUT#9	IN#1	1.35553E-19
C174	IN#1	OUT#2	1.50643E-19
C175	IN#10	OUT#4	1.53813E-19
C176	IN#11	OUT#2	1.59468E-19
C177	OUT#9	IN#8	1.71892E-19
C178	IN#3	OUT#1	1.96134E-19
C179	IN#1	OUT#10	2.05294E-19
C180	OUT#5	IN#7	2.21273E-19
C181	IN	OUT#1	2.30506E-19
C182	OUT#3	IN#11	2.32306E-19
C183	OUT	IN#6	2.68416E-19
C184	IN#3	OUT#10	2.86458E-19
C185	IN#5	OUT#8	3.11517E-19
C186	IN#4	OUT#2	3.39002E-19
C187	OUT#6	IN#9	3.75363E-19
C188	IN#10	OUT#2	4.00049E-19
C189	IN#4	OUT#8	4.11199E-19
C190	IN#1	OUT#1	4.49144E-19
C191	IN#7	OUT#2	4.82054E-19
C192	OUT#3	IN#3	5.28789E-19
C193	IN#10	OUT#3	6.13098E-19
C194	OUT#6	IN#8	6.23542E-19
C195	OUT#9	IN#3	6.31973E-19
C196	OUT#6	IN#6	6.64643E-19
C197	IN#1	OUT#3	6.7634E-19
C198	OUT#3	IN#7	7.58309E-19
C199	OUT#4	IN#7	7.73933E-19
C200	IN#4	OUT#3	8.81042E-19
C201	IN#9	OUT#10	9.05795E-19
C202	OUT#4	IN#3	1.01067E-18
C203	OUT	IN#4	1.10528E-18
C204	VDD#5	VSS#2	6.80575E-20
C205	VSS#3	VDD#5	7.28626E-20
C206	VSS#3	VDD#6	8.04391E-20
C207	VSS#1	VDD#6	1.09976E-19
C208	VDD#2	VSS#2	1.24488E-19
C209	VDD	VSS#3	1.42493E-19
C210	VSS#3	IN#4	6.14226E-20
C211	VSS#1	IN#7	9.21184E-20
C212	IN#5	VSS#2	9.69757E-20
C213	IN#4	VSS#2	1.20518E-19
C214	VSS#3	IN#1	1.68926E-19
C215	VSS#3	IN#8	1.82454E-19
C216	VDD#1	IN#9	1.69709E-19
C217	IN#10	VDD#1	1.87336E-19
C218	VDD#3	IN#6	2.00911E-19
C219	VDD#4	IN#7	2.2286E-19
C220	IN#10	VDD#4	2.29256E-19
C221	VDD	IN#9	2.3727E-19
C222	VDD#5	IN#7	2.47115E-19
C223	VDD	IN#5	2.61028E-19
C224	VDD	IN#4	2.75625E-19
C225	VDD#1	IN#8	2.78472E-19
C226	VDD	IN#1	3.74293E-19
C227	IN	VDD#6	3.84157E-19
C228	IN	VDD#5	4.08364E-19
C229	VDD#3	IN#9	4.45795E-19
C230	VDD	IN#3	5.89631E-19
C231	IN#5	VDD#3	6.28412E-19
C232	IN#3	VDD#6	6.34168E-19
C233	VDD	IN#8	6.63471E-19
C234	VDD#1	IN#6	6.9583E-19
C235	IN#3	VDD#5	7.78185E-19
C236	VDD#2	IN#6	7.94237E-19
C237	IN#4	VDD#3	8.04606E-19
C238	VDD#4	IN#3	8.11498E-19
C239	IN#1	VDD#6	9.94192E-19
C240	IN#1	VDD#5	1.06239E-18
C241	OUT	VSS	6.1205E-17
C242	VDD	VSS	3.38905E-17
C243	IN	VSS	8.26837E-17
C244	IN#10	VSS	4.0838E-17
C245	OUT#9	VSS	1.84609E-18
C246	OUT#6	VSS	5.64525E-17
C247	VDD#1	VSS	7.19481E-17
C248	OUT#5	VSS	3.02749E-17
C249	IN#1	VSS	3.53395E-17
C250	VDD#2	VSS	4.29216E-17
C251	OUT#4	VSS	3.59463E-17
C252	IN#4	VSS	4.34823E-17
C253	VDD#4	VSS	4.07361E-17
C254	OUT#3	VSS	5.05705E-17
C255	IN#5	VSS	9.7473E-17
C256	VDD#5	VSS	1.109E-16
C257	IN#3	VSS	3.59339E-17
C258	VDD#3	VSS	9.39719E-17
C259	IN#6	VSS	6.45259E-17
C260	OUT#8	VSS	2.0916E-17
C261	IN#8	VSS	1.38517E-17
C262	OUT#1	VSS	2.53289E-17
C263	VDD#6	VSS	4.10151E-17
C264	IN#7	VSS	4.67281E-18
C265	IN#9	VSS	6.23512E-18
C266	IN#11	VSS	1.18821E-17
C267	OUT#2	VSS	6.96803E-18
C268	OUT#10	VSS	5.98193E-18
*
*
.ENDS S3D_inv
*
