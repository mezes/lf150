*
*
*
*                       LINUX           Sat Mar 19 18:34:20 2016
*
*
*
*  PROGRAM  advgen
*
*  Name           : advgen - Quantus QRC - (64-bit)
*  Version        : 14.2.3-s099
*  Build Date     : Wed Jun 17 00:01:02 PDT 2015
*
*  HSPICE LIBRARY
*
*
*
*
.SUBCKT test_rppoly A D C
*
*
*  caps2d version: 10
*
*
*       CANONICAL RESISTOR AND CAP/DIODE CARDS
*
RI0	C#4	A#2	resistor 	 6710.0000	L=0.00002U	W=0U
+ $SUB=D#1 
*
*       PARASITIC RESISTOR AND CAP/DIODE CARDS
*
Rm1	A#1	A#2	    1.1800	$L=0.59U	$W=5U
Rm2	C#4	C#2	    2.1800	$L=0.59U	$W=5U
Rl1	A	A#1	    1.0943	$L=1.96U	$W=4.99U
Rl2	C#1	C#2	2.688E-02	$L=0.56U	$W=5U
Rl3	C	C#3	2.688E-02	$L=0.56U	$W=5U
Rl4	C#1	C#3	    0.1578	$L=1.1705U	$W=1.78U
Rl5	D	D#1	    0.4363	$L=3.49U	$W=1.92U
*
*       CAPACITOR CARDS
*
*
C1	A	X3/4	2.83994E-17
C2	A	X3/5	2.74758E-17
C3	X3/4	X3/5	4.25276E-17
C4	X3/4	A#2	3.47804E-17
C5	X3/4	C#4	3.35445E-17
C6	X3/4	A#1	1.01545E-16
C7	X3/4	C#2	2.79076E-17
C8	X3/4	C#1	8.08399E-17
C9	X3/4	C#3	9.77956E-18
C10	X3/5	A#2	3.54914E-17
C11	X3/5	C#4	3.28912E-17
C12	X3/5	A#1	1.06094E-16
C13	X3/5	C#2	2.81585E-17
C14	X3/5	C#1	1.66346E-17
C15	X3/5	C#3	7.33183E-17
C16	A	D	6.66304E-16
C17	X3/4	D	1.16873E-14
C18	X3/5	D	1.17339E-14
C19	A#2	D	3.74859E-16
C20	C#4	D	3.54545E-16
C21	A#1	D	7.36418E-16
C22	C#2	D	4.46936E-16
C23	C#1	D	4.15237E-16
C24	C#3	D	2.85146E-16
*
*
.ENDS test_rppoly
*
